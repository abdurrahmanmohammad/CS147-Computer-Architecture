`timescale 1ns/1ps
module barrel_shifter_tb;
reg [31:0] operand;
reg [31:0] shift;
reg leftNotRight;
wire [31:0] result;
SHIFT32 shifter_inst(.Y(result), .D(operand), .S(shift), .LnR(leftNotRight));
initial begin
	#5;
	#5 operand='b1; shift='b1; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b10000000000000000000000000000000; shift='b1; leftNotRight='b0;
	#5 golden(result,'b1000000000000000000000000000000, operand, shift, leftNotRight);
	#5 operand='b10; shift='b10; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b100; shift='b10; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b100; shift='b11; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b11000; shift='b11; leftNotRight='b0;
	#5 golden(result,'b11, operand, shift, leftNotRight);
	#5 operand='b10000000000000000000000000000000; shift='b1; leftNotRight='b0;
	#5 golden(result,'b1000000000000000000000000000000, operand, shift, leftNotRight);
	#5 operand='b1; shift='b101; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b10000000000000000000000000000000; shift='b1; leftNotRight='b0;
	#5 golden(result,'b1000000000000000000000000000000, operand, shift, leftNotRight);
	#5 operand='b10; shift='b10000; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b100; shift='b10; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b100; shift='b11; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b11000; shift='b11; leftNotRight='b0;
	#5 golden(result,'b11, operand, shift, leftNotRight);
	#5 operand='b11111111111111111111111111111111; shift='b1; leftNotRight='b0;
	#5 golden(result,'b1111111111111111111111111111111, operand, shift, leftNotRight);
	#5 operand='b11111111111111111111111111111111; shift='b10000; leftNotRight='b0;
	#5 golden(result,'b1111111111111111, operand, shift, leftNotRight);
	#5 operand='b11111111111111111111111111111111; shift='b11111; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b10000000000000000000000000000000; shift='b11111; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b1; shift='b1; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b10; shift='b1; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b11; shift='b1; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b100; shift='b1; leftNotRight='b0;
	#5 golden(result,'b10, operand, shift, leftNotRight);
	#5 operand='b101; shift='b1; leftNotRight='b0;
	#5 golden(result,'b10, operand, shift, leftNotRight);
	#5 operand='b110; shift='b1; leftNotRight='b0;
	#5 golden(result,'b11, operand, shift, leftNotRight);
	#5 operand='b111; shift='b1; leftNotRight='b0;
	#5 golden(result,'b11, operand, shift, leftNotRight);
	#5 operand='b1001; shift='b1; leftNotRight='b0;
	#5 golden(result,'b100, operand, shift, leftNotRight);
	#5 operand='b1010; shift='b1; leftNotRight='b0;
	#5 golden(result,'b101, operand, shift, leftNotRight);
	#5 operand='b1011; shift='b1; leftNotRight='b0;
	#5 golden(result,'b101, operand, shift, leftNotRight);
	#5 operand='b1100; shift='b1; leftNotRight='b0;
	#5 golden(result,'b110, operand, shift, leftNotRight);
	#5 operand='b1101; shift='b1; leftNotRight='b0;
	#5 golden(result,'b110, operand, shift, leftNotRight);
	#5 operand='b1110; shift='b1; leftNotRight='b0;
	#5 golden(result,'b111, operand, shift, leftNotRight);
	#5 operand='b1111; shift='b1; leftNotRight='b0;
	#5 golden(result,'b111, operand, shift, leftNotRight);
	#5 operand='b0; shift='b10; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b1; shift='b10; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b10; shift='b10; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b11; shift='b10; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b100; shift='b10; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b101; shift='b10; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b110; shift='b10; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b111; shift='b10; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b1001; shift='b10; leftNotRight='b0;
	#5 golden(result,'b10, operand, shift, leftNotRight);
	#5 operand='b1010; shift='b10; leftNotRight='b0;
	#5 golden(result,'b10, operand, shift, leftNotRight);
	#5 operand='b1011; shift='b10; leftNotRight='b0;
	#5 golden(result,'b10, operand, shift, leftNotRight);
	#5 operand='b1100; shift='b10; leftNotRight='b0;
	#5 golden(result,'b11, operand, shift, leftNotRight);
	#5 operand='b1101; shift='b10; leftNotRight='b0;
	#5 golden(result,'b11, operand, shift, leftNotRight);
	#5 operand='b1110; shift='b10; leftNotRight='b0;
	#5 golden(result,'b11, operand, shift, leftNotRight);
	#5 operand='b1111; shift='b10; leftNotRight='b0;
	#5 golden(result,'b11, operand, shift, leftNotRight);
	#5 operand='b0; shift='b11; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b1; shift='b11; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b10; shift='b11; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b11; shift='b11; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b100; shift='b11; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b101; shift='b11; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b110; shift='b11; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b111; shift='b11; leftNotRight='b0;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b1001; shift='b11; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b1010; shift='b11; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b1011; shift='b11; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight); 
	#5 operand='b1100; shift='b11; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b1101; shift='b11; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b1110; shift='b11; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b1111; shift='b11; leftNotRight='b0;
	#5 golden(result,'b1, operand, shift, leftNotRight);
	#5 operand='b1; shift='b1; leftNotRight='b1;
	#5 golden(result,'b10, operand, shift, leftNotRight);
	#5 operand='b10000000000000000000000000000000; shift='b1; leftNotRight='b1;
	#5 golden(result, 'b100000000000000000000000000000000, operand, shift, leftNotRight);
	#5 operand='b10; shift='b10; leftNotRight='b1;
	#5 golden(result,'b1000, operand, shift, leftNotRight);
	#5 operand='b100; shift='b10; leftNotRight='b1;
	#5 golden(result,'b10000, operand, shift, leftNotRight);
	#5 operand='b100; shift='b11; leftNotRight='b1;
	#5 golden(result,'b100000, operand, shift, leftNotRight);
	#5 operand='b11000; shift='b11; leftNotRight='b1;
	#5 golden(result,'b11000000, operand, shift, leftNotRight);
	#5 operand='b10000000000000000000000000000000; shift='b1; leftNotRight='b1;
	#5 golden(result,'b100000000000000000000000000000000, operand, shift, leftNotRight);
	#5 operand='b1; shift='b101; leftNotRight='b1;
	#5 golden(result,'b100000, operand, shift, leftNotRight);
	#5 operand='b10000000000000000000000000000000; shift='b1; leftNotRight='b1;
	#5 golden(result,'b100000000000000000000000000000000, operand, shift, leftNotRight);
	#5 operand='b10; shift='b10000; leftNotRight='b1;
	#5 golden(result,'b100000000000000000, operand, shift, leftNotRight);
	#5 operand='b100; shift='b10; leftNotRight='b1;
	#5 golden(result,'b10000, operand, shift, leftNotRight);
	#5 operand='b100; shift='b11; leftNotRight='b1;
	#5 golden(result,'b100000, operand, shift, leftNotRight);
	#5 operand='b11111111111111000; shift='b10000; leftNotRight='b1;
	#5 golden(result,'b111111111111110000000000000000000, operand, shift, leftNotRight);
	#5 operand='b11111111111111111111111111111111 ; shift='b1; leftNotRight='b1;
	#5 golden(result,'b11111111111111111111111111111110, operand, shift, leftNotRight);
	#5 operand='b11111111111111111111111111111111; shift='b10; leftNotRight='b1;
	#5 golden(result,'b11111111111111111111111111111100, operand, shift, leftNotRight);
	#5 operand='b11111111111111111111111111111111; shift='b11111; leftNotRight='b1;
	#5 golden(result,'b10000000000000000000000000000000, operand, shift, leftNotRight);
	#5 operand='b10000000000000000000000000000000; shift='b11111; leftNotRight='b1;
	#5 golden(result,'b0, operand, shift, leftNotRight);
	#5 operand='b10000000000000000000000000000000; shift='b1; leftNotRight='b1;
	#5 golden(result,'b0, operand, shift, leftNotRight);
end
task golden;
input [31:0] calculated;
input [31:0] expected;
input [31:0] operand;
input [31:0] shift;
input leftNotRight; 
begin
$write("%d << %d = %d ==> got %d", operand, shift, expected, calculated);
if (calculated == expected) begin
	$write("[PASSED]");
end else if(leftNotRight) begin
	$write("[FAILED]");
end else begin
	$write("[FAILED]");
end
$write("\nRun barrel shift TB\n");
end
endtask
endmodule 